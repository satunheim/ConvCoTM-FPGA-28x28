test 2.vhd here we can ...
